module main;
  initial 
    begin
      $display("Hello world!");
      $finish;
    end
endmodule

// from http://en.wikipedia.org/wiki/Verilog#Example
// Text is available under the Creative Commons Attribution-ShareAlike License
