
class someclass;

  extern function void
    something();

endclass : someclass

