
`include "test.svh"

function void
  someclass::something();

  $display("Something called!");

endfunction : something

